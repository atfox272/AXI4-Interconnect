module sa_RDATA_channel 
#(

)
(
);

endmodule